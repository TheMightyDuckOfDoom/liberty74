VERSION 5.7 ;
BUSBITCHARS "<>" ;
DIVIDERCHAR "/" ;

SITE CoreSite
  CLASS CORE ;
  SYMMETRY R90 ;
  SIZE 0.1 BY 3.6 ;
END CoreSite

MACRO BUF_74LVC1G125
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 3.0 BY 3.6 ;
  SYMMETRY R90 ;
  SITE CoreSite ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
    END
  END A
END BUF_74LVC1G125

MACRO INV_74LVC1G04
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 3.0 BY 3.6 ;
  SYMMETRY R90 ;
  SITE CoreSite ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
    END
  END A
END INV_74LVC1G04

MACRO NAND2_74LVC1G00
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 3.0 BY 3.6 ;
  SYMMETRY R90 ;
  SITE CoreSite ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
    END
  END B
END NAND2_74LVC1G00

MACRO DFFR_74LVC1G175
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 3.0 BY 3.6 ;
  SYMMETRY R90 ;
  SITE CoreSite ;

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
    END
  END D
  PIN RST_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
    END
  END RST_N
END DFFR_74LVC1G175

