VERSION 5.7 ;
BUSBITCHARS "<>" ;
DIVIDERCHAR "/" ;

SITE CoreSite
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.5 BY 3.6 ;
END CoreSite

MACRO BUF_74LVC1G125
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 3.5 BY 3.6 ;
  SYMMETRY R90 ;
  SITE CoreSite ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.25 1.515 0.95 2.025 ;
      LAYER Metal2 ;
        RECT 0.25 1.515 0.95 2.025 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.57 0.565 3.27 1.075 ;
      LAYER Metal2 ;
        RECT 2.57 0.565 3.27 1.075 ;
    END
  END Y
END BUF_74LVC1G125

MACRO NOT_74LVC1G04
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 3.5 BY 3.6 ;
  SYMMETRY R90 ;
  SITE CoreSite ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.25 1.515 0.95 2.025 ;
      LAYER Metal2 ;
        RECT 0.25 1.515 0.95 2.025 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.57 0.565 3.27 1.075 ;
      LAYER Metal2 ;
        RECT 2.57 0.565 3.27 1.075 ;
    END
  END Y
END NOT_74LVC1G04

MACRO AND_74LVC1G08
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 3.5 BY 3.6 ;
  SYMMETRY R90 ;
  SITE CoreSite ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.25 2.465 0.95 2.975 ;
      LAYER Metal2 ;
        RECT 0.25 2.465 0.95 2.975 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.25 1.515 0.95 2.025 ;
      LAYER Metal2 ;
        RECT 0.25 1.515 0.95 2.025 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.57 0.565 3.27 1.075 ;
      LAYER Metal2 ;
        RECT 2.57 0.565 3.27 1.075 ;
    END
  END Y
END AND_74LVC1G08

MACRO NAND_74LVC1G00
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 3.5 BY 3.6 ;
  SYMMETRY R90 ;
  SITE CoreSite ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.25 2.465 0.95 2.975 ;
      LAYER Metal2 ;
        RECT 0.25 2.465 0.95 2.975 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.25 1.515 0.95 2.025 ;
      LAYER Metal2 ;
        RECT 0.25 1.515 0.95 2.025 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.57 0.565 3.27 1.075 ;
      LAYER Metal2 ;
        RECT 2.57 0.565 3.27 1.075 ;
    END
  END Y
END NAND_74LVC1G00

MACRO NOR_74LVC1G02
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 3.5 BY 3.6 ;
  SYMMETRY R90 ;
  SITE CoreSite ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.25 2.465 0.95 2.975 ;
      LAYER Metal2 ;
        RECT 0.25 2.465 0.95 2.975 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.25 1.515 0.95 2.025 ;
      LAYER Metal2 ;
        RECT 0.25 1.515 0.95 2.025 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.57 0.565 3.27 1.075 ;
      LAYER Metal2 ;
        RECT 2.57 0.565 3.27 1.075 ;
    END
  END Y
END NOR_74LVC1G02

MACRO OR_74LVC1G32
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 3.5 BY 3.6 ;
  SYMMETRY R90 ;
  SITE CoreSite ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.25 2.465 0.95 2.975 ;
      LAYER Metal2 ;
        RECT 0.25 2.465 0.95 2.975 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.25 1.515 0.95 2.025 ;
      LAYER Metal2 ;
        RECT 0.25 1.515 0.95 2.025 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.57 0.565 3.27 1.075 ;
      LAYER Metal2 ;
        RECT 2.57 0.565 3.27 1.075 ;
    END
  END Y
END OR_74LVC1G32

MACRO XOR_74LVC1G86
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 3.5 BY 3.6 ;
  SYMMETRY R90 ;
  SITE CoreSite ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.25 2.465 0.95 2.975 ;
      LAYER Metal2 ;
        RECT 0.25 2.465 0.95 2.975 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.25 1.515 0.95 2.025 ;
      LAYER Metal2 ;
        RECT 0.25 1.515 0.95 2.025 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.57 0.565 3.27 1.075 ;
      LAYER Metal2 ;
        RECT 2.57 0.565 3.27 1.075 ;
    END
  END Y
END XOR_74LVC1G86

MACRO DFFSR_74LVC1G74
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 5.9 BY 3.6 ;
  SYMMETRY R90 ;
  SITE CoreSite ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.25 1.895 1.35 2.295 ;
      LAYER Metal2 ;
        RECT 0.25 1.895 1.35 2.295 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.25 2.545 1.35 2.945 ;
      LAYER Metal2 ;
        RECT 0.25 2.545 1.35 2.945 ;
    END
  END C
  PIN RDN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.55 1.245 5.65 1.645 ;
      LAYER Metal2 ;
        RECT 4.55 1.245 5.65 1.645 ;
    END
  END RDN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.55 0.595 5.65 0.995 ;
      LAYER Metal2 ;
        RECT 4.55 0.595 5.65 0.995 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.25 1.245 1.35 1.645 ;
      LAYER Metal2 ;
        RECT 0.25 1.245 1.35 1.645 ;
    END
  END QN
END DFFSR_74LVC1G74