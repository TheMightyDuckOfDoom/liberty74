module \$_NOT_ (input A, output Y);
  \$_NAND_ _TECHMAP_REPLACE_ (.A(A), .B(A), .Y(Y));
endmodule