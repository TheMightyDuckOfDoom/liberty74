VERSION 5.7 ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

PROPERTYDEFINITIONS
  LAYER routingPitch REAL ;
  LAYER routingGrid REAL ;
END PROPERTYDEFINITIONS

LAYER Metal1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.3 ;
  WIDTH 0.13 ;
  SPACING 0.13 ;
end Metal1

LAYER Via1
  TYPE CUT ;
  SPACING 0.5 ;
  WIDTH 0.4 ;
  ENCLOSURE 0.13 0.13 ;
END Via1

LAYER Metal2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.3 ;
  WIDTH 0.13 ;
  SPACING 0.13 ;
end Metal2

VIA Via1_0 DEFAULT
  LAYER Metal1 ;
    RECT -0.33 -0.33 0.33 0.33 ;
  LAYER Via1 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER Metal2 ;
    RECT -0.33 -0.33 0.33 0.33 ;
END Via1_0
